library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package	constants is
        type TPicoType is ( pbtI, pbtII, pbt3, pbtS ) ;
	constant PicoType : TPicoType := pbt3 ;
	CONSTANT ADDRSIZE : natural := 10;
	CONSTANT INSTSIZE : natural := 18;
	CONSTANT JADDRSIZE : natural := 11;
	CONSTANT JDATASIZE : natural := 9;
end package ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

library unisim ;
use unisim.vcomponents.all ;

use work.constants.all;

entity prog_rom is
    port ( 
        clk : in std_logic ;
        reset : out std_logic ;
        address : in std_logic_vector( ADDRSIZE - 1 downto 0 ) ;
        instruction : out std_logic_vector( INSTSIZE - 1 downto 0 )
    ) ;
end entity prog_rom ;

architecture mix of prog_rom is
    component jtag_shifter is
        port ( 
			clk : in std_logic ;
			user1 : out std_logic ;
            write : out std_logic ;
            addr : out std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
            data : out std_logic_vector( JDATASIZE - 1 downto 0 )
        ) ;
    end component ;

    signal jaddr : std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
    signal jdata : std_logic_vector( JDATASIZE - 1 downto 0 ) ;
    signal juser1 : std_logic ;
    signal jwrite : std_logic ;

    attribute INIT_00 : string ;
    attribute INIT_01 : string ;
    attribute INIT_02 : string ;
    attribute INIT_03 : string ;
    attribute INIT_04 : string ;
    attribute INIT_05 : string ;
    attribute INIT_06 : string ;
    attribute INIT_07 : string ;
    attribute INIT_08 : string ;
    attribute INIT_09 : string ;
    attribute INIT_0A : string ;
    attribute INIT_0B : string ;
    attribute INIT_0C : string ;
    attribute INIT_0D : string ;
    attribute INIT_0E : string ;
    attribute INIT_0F : string ;
    attribute INIT_10 : string ;
    attribute INIT_11 : string ;
    attribute INIT_12 : string ;
    attribute INIT_13 : string ;
    attribute INIT_14 : string ;
    attribute INIT_15 : string ;
    attribute INIT_16 : string ;
    attribute INIT_17 : string ;
    attribute INIT_18 : string ;
    attribute INIT_19 : string ;
    attribute INIT_1A : string ;
    attribute INIT_1B : string ;
    attribute INIT_1C : string ;
    attribute INIT_1D : string ;
    attribute INIT_1E : string ;
    attribute INIT_1F : string ;
    attribute INIT_20 : string ;
    attribute INIT_21 : string ;
    attribute INIT_22 : string ;
    attribute INIT_23 : string ;
    attribute INIT_24 : string ;
    attribute INIT_25 : string ;
    attribute INIT_26 : string ;
    attribute INIT_27 : string ;
    attribute INIT_28 : string ;
    attribute INIT_29 : string ;
    attribute INIT_2A : string ;
    attribute INIT_2B : string ;
    attribute INIT_2C : string ;
    attribute INIT_2D : string ;
    attribute INIT_2E : string ;
    attribute INIT_2F : string ;
    attribute INIT_30 : string ;
    attribute INIT_31 : string ;
    attribute INIT_32 : string ;
    attribute INIT_33 : string ;
    attribute INIT_34 : string ;
    attribute INIT_35 : string ;
    attribute INIT_36 : string ;
    attribute INIT_37 : string ;
    attribute INIT_38 : string ;
    attribute INIT_39 : string ;
    attribute INIT_3A : string ;
    attribute INIT_3B : string ;
    attribute INIT_3C : string ;
    attribute INIT_3D : string ;
    attribute INIT_3E : string ;
    attribute INIT_3F : string ;
    attribute INITP_00 : string ;
    attribute INITP_01 : string ;
    attribute INITP_02 : string ;
    attribute INITP_03 : string ;
    attribute INITP_04 : string ;
    attribute INITP_05 : string ;
    attribute INITP_06 : string ;
    attribute INITP_07 : string ;
begin
	I18: IF PicoType = pbt3 GENERATE
  	    attribute INIT_00 of bram : label is "400040C001105C09EF00CE01009E0EF40F0100580106052000120106051000F0" ;
	    attribute INIT_01 of bram : label is "00C6054200C6055200C6054900C6054500C6055300C6054E00C6054540075513" ;
	    attribute INIT_02 of bram : label is "00C6056300C6056500C6057600C60561009200C6054400C6054300C6054C0092" ;
	    attribute INIT_03 of bram : label is "056500C6057200C6057200C605450101A00000C6054D00C6054F00C605520092" ;
	    attribute INIT_04 of bram : label is "413600C605320038413600C605310038A00000C6052000C6057200C6057500C6" ;
	    attribute INIT_05 of bram : label is "00C6056D00C6056D00C6056F00C60543413600C605300038413600C605330038" ;
	    attribute INIT_06 of bram : label is "00C60573009200C6056E00C60575009200C6057200C6056500C6057400C60575" ;
	    attribute INIT_07 of bram : label is "057400C6056500C60528009200C6056800C6056300C6057400C6056900C60577" ;
	    attribute INIT_08 of bram : label is "052900C6056C00C6057500C6056500C60573009200C6056E00C60575009200C6" ;
	    attribute INIT_09 of bram : label is "00990219A000549AC10100950128A0005496C001000BA00000C60520A00000C6" ;
	    attribute INIT_0A of bram : label is "0095C4A0E401A00054A9C40100A30432A00054A4C301009E0314A000549FC201" ;
	    attribute INIT_0B of bram : label is "0406040604071450009500B3C408A4F01450A00000ADC4A0A4F8A000C4A0E401" ;
	    attribute INIT_0C of bram : label is "0406040704071450009500ADC4A0C40CA4F01450A000C4A004F0009900B30406" ;
	    attribute INIT_0D of bram : label is "0095C4A0E40145800095C4A0E401C4A0040EA000C4A004F0009900ADC4A00406" ;
	    attribute INIT_0E of bram : label is "A0000099C4A00404D500000E000E000E000EA5F0C4A0E40140800095C4A0E401" ;
	    attribute INIT_0F of bram : label is "050C00B7050600B70528009900B30420009900B3009E00B300A300B3043000A3" ;
	    attribute INIT_10 of bram : label is "A00000B7C5C0A50FA00000B7C580A50F510C2510A000009E009E00B7050100B7" ;
	    attribute INIT_11 of bram : label is "8301938058305123C0018301504C49005930512F400040C00300A00000B70518" ;
	    attribute INIT_12 of bram : label is "41C04127513AC701512FC801830100C655300710830158300101411B504CC901" ;
	    attribute INIT_13 of bram : label is "00000000412707C801060520A0000106051041364113512F40005130501040C0" ;
	    attribute INIT_14 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_15 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_16 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_17 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_18 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_19 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_20 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_21 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_22 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_23 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_24 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_25 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_26 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_27 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_28 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_29 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_30 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_31 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_32 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_33 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_34 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_35 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_36 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_37 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_38 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_39 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_00 of bram : label is "333CCCCCCF33CCCCCCCCF3F3F3F3B3333333B333CCCCF333CCCCCCCF4F5C3CF3" ;
	    attribute INITP_01 of bram : label is "333CFFF3B82A8838E0E228FAA8F80A3EA8F02E28E2DCB72DCB72D2CB33333CCF" ;
	    attribute INITP_02 of bram : label is "000000000000000000000000000000000CCB3F743DD704FD535D342CB0B0DBF3" ;
	    attribute INITP_03 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_07 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
	            INIT_00 => X"400040C001105C09EF00CE01009E0EF40F0100580106052000120106051000F0",
	            INIT_01 => X"00C6054200C6055200C6054900C6054500C6055300C6054E00C6054540075513",
	            INIT_02 => X"00C6056300C6056500C6057600C60561009200C6054400C6054300C6054C0092",
	            INIT_03 => X"056500C6057200C6057200C605450101A00000C6054D00C6054F00C605520092",
	            INIT_04 => X"413600C605320038413600C605310038A00000C6052000C6057200C6057500C6",
	            INIT_05 => X"00C6056D00C6056D00C6056F00C60543413600C605300038413600C605330038",
	            INIT_06 => X"00C60573009200C6056E00C60575009200C6057200C6056500C6057400C60575",
	            INIT_07 => X"057400C6056500C60528009200C6056800C6056300C6057400C6056900C60577",
	            INIT_08 => X"052900C6056C00C6057500C6056500C60573009200C6056E00C60575009200C6",
	            INIT_09 => X"00990219A000549AC10100950128A0005496C001000BA00000C60520A00000C6",
	            INIT_0A => X"0095C4A0E401A00054A9C40100A30432A00054A4C301009E0314A000549FC201",
	            INIT_0B => X"0406040604071450009500B3C408A4F01450A00000ADC4A0A4F8A000C4A0E401",
	            INIT_0C => X"0406040704071450009500ADC4A0C40CA4F01450A000C4A004F0009900B30406",
	            INIT_0D => X"0095C4A0E40145800095C4A0E401C4A0040EA000C4A004F0009900ADC4A00406",
	            INIT_0E => X"A0000099C4A00404D500000E000E000E000EA5F0C4A0E40140800095C4A0E401",
	            INIT_0F => X"050C00B7050600B70528009900B30420009900B3009E00B300A300B3043000A3",
	            INIT_10 => X"A00000B7C5C0A50FA00000B7C580A50F510C2510A000009E009E00B7050100B7",
	            INIT_11 => X"8301938058305123C0018301504C49005930512F400040C00300A00000B70518",
	            INIT_12 => X"41C04127513AC701512FC801830100C655300710830158300101411B504CC901",
	            INIT_13 => X"00000000412707C801060520A0000106051041364113512F40005130501040C0",
	            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_00 => X"333CCCCCCF33CCCCCCCCF3F3F3F3B3333333B333CCCCF333CCCCCCCF4F5C3CF3",
	            INITP_01 => X"333CFFF3B82A8838E0E228FAA8F80A3EA8F02E28E2DCB72DCB72D2CB33333CCF",
	            INITP_02 => X"000000000000000000000000000000000CCB3F743DD704FD535D342CB0B0DBF3",
	            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000"
	        )
	        port map (
	            DIB => "0000000000000000",
	            DIPB => "00",
	            ENB => '1',
	            WEB => '0',
	            SSRB => '0',
	            CLKB => clk,
	            ADDRB => address,
	            DOB => instruction( INSTSIZE - 3 downto 0 ),
	            DOPB => instruction( INSTSIZE - 1 downto INSTSIZE - 2 ),
	            DIA => jdata( JDATASIZE - 2 downto 0 ),
	            DIPA => jdata( JDATASIZE - 1 downto JDATASIZE - 1 ),
	            ENA => juser1,
	            WEA => jwrite,
	            SSRA => '0',
	            CLKA => clk,
	            ADDRA => jaddr,
	            DOA => open,
	            DOPA => open 
	        ) ;
	end generate ;

	jdata <= ( others => '0' ) ;
	jaddr <= ( others => '0' ) ;
	juser1 <= '0' ;
	jwrite <= '0' ;
end architecture mix ;
